

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO ULA_com_registrador 
  PIN clk 
    ANTENNAPARTIALMETALAREA 23.492 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.16892 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 45.12 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.7842 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0466374 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.17078 LAYER V3 ;
  END clk
  PIN rst 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.011 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.14 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.2457 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.141714 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.12 LAYER V3 ;
  END rst
  PIN A[31] 
    ANTENNAPARTIALMETALAREA 2.0104 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01436 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 15.9152 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.11424 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.68 LAYER M4 ; 
    ANTENNAMAXAREACAR 28.6 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.208294 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.345882 LAYER V4 ;
  END A[31]
  PIN A[30] 
    ANTENNAPARTIALMETALAREA 0.168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0012 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 4.6256 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0336 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.18 LAYER M4 ; 
    ANTENNAMAXAREACAR 7.53099 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0583071 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.249344 LAYER V4 ;
  END A[30]
  PIN A[29] 
    ANTENNAPARTIALMETALAREA 4.9896 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03564 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 9.016 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06496 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.48 LAYER M4 ; 
    ANTENNAMAXAREACAR 5.17488 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0387744 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.20872 LAYER V4 ;
  END A[29]
  PIN A[28] 
    ANTENNAPARTIALMETALAREA 6.1656 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0446 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.12 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.6692 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0801923 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.297722 LAYER V3 ;
  END A[28]
  PIN A[27] 
    ANTENNAPARTIALMETALAREA 3.108 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.63 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.30554 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0425856 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.293639 LAYER V3 ;
  END A[27]
  PIN A[26] 
    ANTENNAPARTIALMETALAREA 3.6568 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02668 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.3 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.19881 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0326792 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.147925 LAYER V3 ;
  END A[26]
  PIN A[25] 
    ANTENNAPARTIALMETALAREA 12.9864 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09276 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.12 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.54411 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0562385 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.230588 LAYER V3 ;
  END A[25]
  PIN A[24] 
    ANTENNAPARTIALMETALAREA 14.1624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10172 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.28906 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0471165 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.198481 LAYER V3 ;
  END A[24]
  PIN A[23] 
    ANTENNAPARTIALMETALAREA 7.3416 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05244 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 6.1936 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0448 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 6.14738 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0465051 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.215712 LAYER V4 ;
  END A[23]
  PIN A[22] 
    ANTENNAPARTIALMETALAREA 20.4344 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14652 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.07225 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0601434 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.230588 LAYER V3 ;
  END A[22]
  PIN A[21] 
    ANTENNAPARTIALMETALAREA 16.2792 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.11628 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.92138 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0436756 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.147925 LAYER V3 ;
  END A[21]
  PIN A[20] 
    ANTENNAPARTIALMETALAREA 15.3384 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.67331 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0669363 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.254346 LAYER V3 ;
  END A[20]
  PIN A[19] 
    ANTENNAPARTIALMETALAREA 13.6136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09724 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.2 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.90952 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0509746 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0926289 LAYER V3 ;
  END A[19]
  PIN A[18] 
    ANTENNAPARTIALMETALAREA 19.7288 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14092 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.87 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.31018 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0600958 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.122077 LAYER V3 ;
  END A[18]
  PIN A[17] 
    ANTENNAPARTIALMETALAREA 17.3768 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.12412 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 10.2704 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.07392 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.63 LAYER M4 ; 
    ANTENNAMAXAREACAR 5.95183 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.045869 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.201404 LAYER V4 ;
  END A[17]
  PIN A[16] 
    ANTENNAPARTIALMETALAREA 28.9016 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.207 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.3 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.29068 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.060224 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0887547 LAYER V3 ;
  END A[16]
  PIN A[15] 
    ANTENNAPARTIALMETALAREA 34.86 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.24956 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.8241 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0795237 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.203636 LAYER V3 ;
  END A[15]
  PIN A[14] 
    ANTENNAPARTIALMETALAREA 0.4424 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00316 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 4.9392 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03584 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 12.8921 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0969403 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.149756 LAYER V4 ;
  END A[14]
  PIN A[13] 
    ANTENNAPARTIALMETALAREA 33.684 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2406 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.52 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.1738 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0805035 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.129587 LAYER V3 ;
  END A[13]
  PIN A[12] 
    ANTENNAPARTIALMETALAREA 31.0184 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22156 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.0643 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0741864 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.198481 LAYER V3 ;
  END A[12]
  PIN A[11] 
    ANTENNAPARTIALMETALAREA 1.6968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01212 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.176 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00896 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 10.8798 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0801005 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.314952 LAYER V4 ;
  END A[11]
  PIN A[10] 
    ANTENNAPARTIALMETALAREA 3.5784 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.02556 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 1.4896 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0112 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 8.01824 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0590194 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.133702 LAYER V4 ;
  END A[10]
  PIN A[9] 
    ANTENNAPARTIALMETALAREA 6.4008 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04572 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 12.3088 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.08848 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.24 LAYER M4 ; 
    ANTENNAMAXAREACAR 9.46396 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0695547 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.288835 LAYER V4 ;
  END A[9]
  PIN A[8] 
    ANTENNAPARTIALMETALAREA 12.9864 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09276 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 6.664 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04816 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 9.20185 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0683333 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.159902 LAYER V4 ;
  END A[8]
  PIN A[7] 
    ANTENNAPARTIALMETALAREA 1.2264 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00876 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 8.5456 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0616 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 12.1861 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.089515 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.185858 LAYER V4 ;
  END A[7]
  PIN A[6] 
    ANTENNAPARTIALMETALAREA 2.324 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0166 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 11.368 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.08176 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 13.4706 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0993371 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.247819 LAYER V4 ;
  END A[6]
  PIN A[5] 
    ANTENNAPARTIALMETALAREA 1.6968 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01212 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.3136 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0028 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V4 ;
    ANTENNAPARTIALMETALAREA 38.4944 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 0.27552 LAYER MT ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER MT ; 
    ANTENNAMAXAREACAR 14.483 LAYER MT ;
    ANTENNAMAXSIDEAREACAR 0.10709 LAYER MT ;
    ANTENNAMAXCUTCAR 0.232943 LAYER FT ;
  END A[5]
  PIN A[4] 
    ANTENNAPARTIALMETALAREA 3.108 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0222 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 7.1344 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05152 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V4 ;
    ANTENNAPARTIALMETALAREA 40.5328 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 0.29008 LAYER MT ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER MT ; 
    ANTENNAMAXAREACAR 12.9239 LAYER MT ;
    ANTENNAMAXSIDEAREACAR 0.095338 LAYER MT ;
    ANTENNAMAXCUTCAR 0.238098 LAYER FT ;
  END A[4]
  PIN A[3] 
    ANTENNAPARTIALMETALAREA 44.0328 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.31452 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.63 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.7801 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0938712 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.132227 LAYER V3 ;
  END A[3]
  PIN A[2] 
    ANTENNAPARTIALMETALAREA 49.2856 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3526 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.3146 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.105079 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.305455 LAYER V3 ;
  END A[2]
  PIN A[1] 
    ANTENNAPARTIALMETALAREA 7.812 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0558 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.392 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00336 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V4 ;
    ANTENNAPARTIALMETALAREA 30.3408 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 0.21728 LAYER MT ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER MT ; 
    ANTENNAMAXAREACAR 12.2828 LAYER MT ;
    ANTENNAMAXSIDEAREACAR 0.0900225 LAYER MT ;
    ANTENNAMAXCUTCAR 0.238098 LAYER FT ;
  END A[1]
  PIN A[0] 
    ANTENNAPARTIALMETALAREA 45.2872 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.32348 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.46 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.5801 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.148381 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.140759 LAYER V3 ;
  END A[0]
  PIN sel[1] 
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.6552 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05468 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.83 LAYER M3 ; 
    ANTENNAMAXAREACAR 4.24933 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0325948 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0856831 LAYER V3 ;
  END sel[1]
  PIN sel[0] 
    ANTENNADIFFAREA 0.16 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 39.6704 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.28672 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 17.05 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.85097 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0737286 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.247008 LAYER V3 ;
  END sel[0]
  PIN S[31] 
    ANTENNAPARTIALMETALAREA 2.0104 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01436 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 0.97 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 2.4304 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01792 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.99 LAYER M4 ; 
    ANTENNAMAXAREACAR 5.08135 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0384702 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.171029 LAYER V4 ;
  END S[31]
  PIN S[30] 
    ANTENNAPARTIALMETALAREA 9.0664 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06476 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.8624 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V4 ;
    ANTENNADIFFAREA 0.97 LAYER MT ; 
    ANTENNAPARTIALMETALAREA 26.1072 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 0.18704 LAYER MT ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.38 LAYER MT ; 
    ANTENNAMAXAREACAR 6.55002 LAYER MT ;
    ANTENNAMAXSIDEAREACAR 0.0492053 LAYER MT ;
    ANTENNAMAXCUTCAR 0.246734 LAYER FT ;
  END S[30]
  PIN S[29] 
    ANTENNAPARTIALMETALAREA 7.4984 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05356 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.3136 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0028 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V4 ;
    ANTENNADIFFAREA 1.62 LAYER MT ; 
    ANTENNAPARTIALMETALAREA 26.5776 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 0.1904 LAYER MT ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER MT ; 
    ANTENNAMAXAREACAR 3.9142 LAYER MT ;
    ANTENNAMAXSIDEAREACAR 0.0297823 LAYER MT ;
    ANTENNAMAXCUTCAR 0.977181 LAYER FT ;
  END S[29]
  PIN S[28] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 47.404 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.33916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.447 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.164524 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.6272 LAYER V3 ;
  END S[28]
  PIN S[27] 
    ANTENNAPARTIALMETALAREA 0.2856 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00204 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 2.5872 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01904 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V4 ;
    ANTENNADIFFAREA 1.62 LAYER MT ; 
    ANTENNAPARTIALMETALAREA 39.7488 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 0.28448 LAYER MT ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.64 LAYER MT ; 
    ANTENNAMAXAREACAR 9.19513 LAYER MT ;
    ANTENNAMAXSIDEAREACAR 0.0682215 LAYER MT ;
    ANTENNAMAXCUTCAR 0.499222 LAYER FT ;
  END S[27]
  PIN S[26] 
    ANTENNAPARTIALMETALAREA 1.0696 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00764 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNAPARTIALMETALAREA 0.8624 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.00672 LAYER M4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V4 ;
    ANTENNADIFFAREA 1.62 LAYER MT ; 
    ANTENNAPARTIALMETALAREA 36.9264 LAYER MT ;
    ANTENNAPARTIALMETALSIDEAREA 0.26432 LAYER MT ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER MT ; 
    ANTENNAMAXAREACAR 9.09936 LAYER MT ;
    ANTENNAMAXSIDEAREACAR 0.0675611 LAYER MT ;
    ANTENNAMAXCUTCAR 0.492526 LAYER FT ;
  END S[26]
  PIN S[25] 
    ANTENNAPARTIALMETALAREA 21.4536 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15324 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 1.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 9.016 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06496 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8 LAYER M4 ; 
    ANTENNAMAXAREACAR 8.95832 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.068232 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.961432 LAYER V4 ;
  END S[25]
  PIN S[24] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 37.1336 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.26636 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.92816 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0302104 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.336259 LAYER V3 ;
  END S[24]
  PIN S[23] 
    ANTENNAPARTIALMETALAREA 3.892 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0278 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 1.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.5072 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04704 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8 LAYER M4 ; 
    ANTENNAMAXAREACAR 3.57616 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.027632 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.354863 LAYER V4 ;
  END S[23]
  PIN S[22] 
    ANTENNAPARTIALMETALAREA 10.7912 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.07708 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 1.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 5.7232 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04144 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M4 ; 
    ANTENNAMAXAREACAR 3.08715 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.024133 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.348062 LAYER V4 ;
  END S[22]
  PIN S[21] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 36.7416 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.263 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.32 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.95018 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.07527 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.6272 LAYER V3 ;
  END S[21]
  PIN S[20] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 35.4088 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.25292 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 14.228 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.105789 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.6272 LAYER V3 ;
  END S[20]
  PIN S[19] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 33.1352 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.23724 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.5 LAYER M3 ; 
    ANTENNAMAXAREACAR 27.2455 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.198808 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.6272 LAYER V3 ;
  END S[19]
  PIN S[18] 
    ANTENNAPARTIALMETALAREA 7.9688 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05692 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 1.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 6.8208 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04928 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 2.66 LAYER M4 ; 
    ANTENNAMAXAREACAR 13.1075 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.107064 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.699989 LAYER V4 ;
  END S[18]
  PIN S[17] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 29.9208 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.21484 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.64 LAYER M3 ; 
    ANTENNAMAXAREACAR 11.3302 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0832522 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.388985 LAYER V3 ;
  END S[17]
  PIN S[16] 
    ANTENNAPARTIALMETALAREA 10.4776 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.07484 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 1.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 8.3888 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.06048 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER M4 ; 
    ANTENNAMAXAREACAR 5.91789 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0481707 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.354449 LAYER V4 ;
  END S[16]
  PIN S[15] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 16.828 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.12076 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.30869 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0614733 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.340176 LAYER V3 ;
  END S[15]
  PIN S[14] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.2408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10172 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 7.60366 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0620358 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.334789 LAYER V3 ;
  END S[14]
  PIN S[13] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 19.2584 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.13868 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.32 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.2978 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0424294 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.9408 LAYER V3 ;
  END S[13]
  PIN S[12] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 22.0808 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.15772 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.87659 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0318499 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.6272 LAYER V3 ;
  END S[12]
  PIN S[11] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 27.02 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.19356 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.3046 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0908562 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.456145 LAYER V3 ;
  END S[11]
  PIN S[10] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 31.6456 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.22716 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.55 LAYER M3 ; 
    ANTENNAMAXAREACAR 20.2099 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.149187 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.9408 LAYER V3 ;
  END S[10]
  PIN S[9] 
    ANTENNAPARTIALMETALAREA 17.6904 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.12636 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 1.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.4688 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03248 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.98 LAYER M4 ; 
    ANTENNAMAXAREACAR 8.06664 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.0618318 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.642943 LAYER V4 ;
  END S[9]
  PIN S[8] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 19.8856 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.14316 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.09546 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0386815 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.40023 LAYER V3 ;
  END S[8]
  PIN S[7] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 17.612 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.12636 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER M3 ; 
    ANTENNAMAXAREACAR 18.3979 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.135601 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.6272 LAYER V3 ;
  END S[7]
  PIN S[6] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.9464 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10732 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.8 LAYER M3 ; 
    ANTENNAMAXAREACAR 10.0616 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.074326 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.456145 LAYER V3 ;
  END S[6]
  PIN S[5] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 14.2408 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.10284 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER M3 ; 
    ANTENNAMAXAREACAR 9.45273 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0717341 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.6272 LAYER V3 ;
  END S[5]
  PIN S[4] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 6.636 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.04796 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.56 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.46649 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0265973 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.384873 LAYER V3 ;
  END S[4]
  PIN S[3] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 8.204 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.05916 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.64 LAYER M3 ; 
    ANTENNAMAXAREACAR 5.51485 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0417147 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.384873 LAYER V3 ;
  END S[3]
  PIN S[2] 
    ANTENNADIFFAREA 1.62 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 15.5736 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1118 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 4.31 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.48592 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0275208 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.9408 LAYER V3 ;
  END S[2]
  PIN S[1] 
    ANTENNAPARTIALMETALAREA 0.168 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0012 LAYER M3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER V3 ;
    ANTENNADIFFAREA 1.62 LAYER M4 ; 
    ANTENNAPARTIALMETALAREA 4.6256 LAYER M4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0336 LAYER M4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.42 LAYER M4 ; 
    ANTENNAMAXAREACAR 33.8466 LAYER M4 ;
    ANTENNAMAXSIDEAREACAR 0.246007 LAYER M4 ;
    ANTENNAMAXCUTCAR 0.650124 LAYER V4 ;
  END S[1]
  PIN S[0] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.7544 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03452 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.87 LAYER M3 ; 
    ANTENNAMAXAREACAR 12.3271 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0942698 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.2455 LAYER V3 ;
  END S[0]
END ULA_com_registrador

END LIBRARY
