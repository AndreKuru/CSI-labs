

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO contador 
  PIN clk 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.011 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.64 LAYER M3 ; 
    ANTENNAMAXAREACAR 3.07333 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0247447 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.0417021 LAYER V3 ;
  END clk
  PIN rst 
    ANTENNAPARTIALMETALAREA 1.8536 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.01324 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.14 LAYER M3 ; 
    ANTENNAMAXAREACAR 22.7257 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.173714 LAYER M3 ;
    ANTENNAMAXCUTCAR 1.12 LAYER V3 ;
  END rst
  PIN count[3] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 4.3624 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.03116 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.77 LAYER M3 ; 
    ANTENNAMAXAREACAR 1.43814 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0122227 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.154716 LAYER V3 ;
  END count[3]
  PIN count[2] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 13.6136 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.09724 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.06 LAYER M3 ; 
    ANTENNAMAXAREACAR 2.64785 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0211881 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.147925 LAYER V3 ;
  END count[2]
  PIN count[1] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 1.54 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.011 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.62 LAYER M3 ; 
    ANTENNAMAXAREACAR 8.22953 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.0700328 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.468395 LAYER V3 ;
  END count[1]
  PIN count[0] 
    ANTENNADIFFAREA 0.97 LAYER M3 ; 
    ANTENNAPARTIALMETALAREA 7.7336 LAYER M3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0558 LAYER M3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.74 LAYER M3 ; 
    ANTENNAMAXAREACAR 6.39428 LAYER M3 ;
    ANTENNAMAXSIDEAREACAR 0.051507 LAYER M3 ;
    ANTENNAMAXCUTCAR 0.423784 LAYER V3 ;
  END count[0]
END contador

END LIBRARY
